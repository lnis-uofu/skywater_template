

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO mips 
  PIN clk 
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.2632 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2932 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 32.564 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 123.575 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 22.1648 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 84.5032 LAYER METAL5 ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 10.3838 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.6069 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 18.872 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 72.0376 LAYER METAL4 ;
  END reset
  PIN memdata[7] 
    ANTENNAPARTIALMETALAREA 5.5734 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0993 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 6.5352 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.0372 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.612 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 40.4708 LAYER METAL4 ;
  END memdata[7]
  PIN memdata[6] 
    ANTENNAPARTIALMETALAREA 14.2534 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 54.5529 LAYER METAL4 ;
  END memdata[6]
  PIN memdata[5] 
    ANTENNAPARTIALMETALAREA 6.9846 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.4417 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.8472 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.158 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.8872 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.9412 LAYER METAL4 ;
  END memdata[5]
  PIN memdata[4] 
    ANTENNAPARTIALMETALAREA 13.6766 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 52.0725 LAYER METAL4 ;
  END memdata[4]
  PIN memdata[3] 
    ANTENNAPARTIALMETALAREA 5.4166 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5057 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.2632 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2932 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 11.0824 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.2516 LAYER METAL4 ;
  END memdata[3]
  PIN memdata[2] 
    ANTENNAPARTIALMETALAREA 0.5558 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1041 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.6152 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1972 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 17.3544 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 65.9956 LAYER METAL4 ;
  END memdata[2]
  PIN memdata[1] 
    ANTENNAPARTIALMETALAREA 4.9462 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.7249 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.5024 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.1384 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 14.4816 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 55.4168 LAYER METAL4 ;
  END memdata[1]
  PIN memdata[0] 
    ANTENNAPARTIALMETALAREA 0.2422 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9169 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 13.8544 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.0424 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 6.5352 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 25.0372 LAYER METAL4 ;
  END memdata[0]
  PIN memread 
    ANTENNAPARTIALMETALAREA 13.2566 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 50.1857 LAYER METAL5 ;
  END memread
  PIN memwrite 
    ANTENNAPARTIALMETALAREA 14.8246 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.1217 LAYER METAL3 ;
  END memwrite
  PIN adr[7] 
    ANTENNAPARTIALMETALAREA 11.0614 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.8753 LAYER METAL3 ;
  END adr[7]
  PIN adr[6] 
    ANTENNAPARTIALMETALAREA 9.6502 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5329 LAYER METAL3 ;
  END adr[6]
  PIN adr[5] 
    ANTENNAPARTIALMETALAREA 12.3158 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.6241 LAYER METAL3 ;
  END adr[5]
  PIN adr[4] 
    ANTENNAPARTIALMETALAREA 8.7094 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.9713 LAYER METAL3 ;
  END adr[4]
  PIN adr[3] 
    ANTENNAPARTIALMETALAREA 11.0614 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.8753 LAYER METAL3 ;
  END adr[3]
  PIN adr[2] 
    ANTENNAPARTIALMETALAREA 11.2182 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.4689 LAYER METAL3 ;
  END adr[2]
  PIN adr[1] 
    ANTENNAPARTIALMETALAREA 9.6502 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.5329 LAYER METAL3 ;
  END adr[1]
  PIN adr[0] 
    ANTENNAPARTIALMETALAREA 9.4934 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 35.9393 LAYER METAL5 ;
  END adr[0]
  PIN writedata[7] 
    ANTENNAPARTIALMETALAREA 0.8694 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.2913 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.42 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8868 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 19.5496 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 74.306 LAYER METAL5 ;
  END writedata[7]
  PIN writedata[6] 
    ANTENNAPARTIALMETALAREA 0.2422 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9169 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.8904 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6676 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 21.588 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 82.0228 LAYER METAL5 ;
  END writedata[6]
  PIN writedata[5] 
    ANTENNAPARTIALMETALAREA 0.7126 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6977 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.7336 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.074 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 20.804 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 79.0548 LAYER METAL5 ;
  END writedata[5]
  PIN writedata[4] 
    ANTENNAPARTIALMETALAREA 25.0166 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 94.7057 LAYER METAL5 ;
  END writedata[4]
  PIN writedata[3] 
    ANTENNAPARTIALMETALAREA 1.183 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4785 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.0472 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.2612 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 26.7624 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 101.612 LAYER METAL4 ;
  END writedata[3]
  PIN writedata[2] 
    ANTENNAPARTIALMETALAREA 33.327 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 126.167 LAYER METAL3 ;
  END writedata[2]
  PIN writedata[1] 
    ANTENNAPARTIALMETALAREA 3.0646 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6017 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.2632 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2932 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 31.416 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 119.526 LAYER METAL5 ;
  END writedata[1]
  PIN writedata[0] 
    ANTENNAPARTIALMETALAREA 33.1198 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 125.679 LAYER METAL3 ;
  END writedata[0]
END mips

END LIBRARY
